`define PRMT 
parameter pckg_sz = 32;
parameter drvrs = 16;
