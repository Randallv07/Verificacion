/*UVM_INFO Driver.sv(59) @ 230: uvm_test_top.amb_inst.agent.drv_inst7 [DRV] Driver #7: Fuente: [4][0], envia el mensaje: 441c al driver destino [3][5], en modo 1
UVM_INFO Driver.sv(59) @ 350: uvm_test_top.amb_inst.agent.drv_inst1 [DRV] Driver #1: Fuente: [0][2], envia el mensaje: 3500 al driver destino [5][2], en modo 0
UVM_INFO Driver.sv(59) @ 510: uvm_test_top.amb_inst.agent.drv_inst15 [DRV] Driver #15: Fuente: [4][5], envia el mensaje: 3a5d al driver destino [4][5], en modo 1
UVM_INFO Driver.sv(59) @ 1350: uvm_test_top.amb_inst.agent.drv_inst5 [DRV] Driver #5: Fuente: [2][0], envia el mensaje: 6fcf al driver destino [1][5], en modo 0
UVM_INFO Driver.sv(59) @ 1450: uvm_test_top.amb_inst.agent.drv_inst3 [DRV] Driver #3: Fuente: [0][4], envia el mensaje: 1154 al driver destino [5][1], en modo 0
UVM_INFO Driver.sv(59) @ 630: uvm_test_top.amb_inst.agent.drv_inst3 [DRV] Driver #3: Fuente: [0][4], envia el mensaje: 1d35 al driver destino [5][3], en modo 1
UVM_INFO Driver.sv(59) @ 770: uvm_test_top.amb_inst.agent.drv_inst6 [DRV] Driver #6: Fuente: [3][0], envia el mensaje: 2a94 al driver destino [5][3], en modo 1
UVM_INFO Driver.sv(59) @ 910: uvm_test_top.amb_inst.agent.drv_inst14 [DRV] Driver #14: Fuente: [3][5], envia el mensaje: 518d al driver destino [5][4], en modo 1
UVM_INFO Driver.sv(59) @ 1010: uvm_test_top.amb_inst.agent.drv_inst1 [DRV] Driver #1: Fuente: [0][2], envia el mensaje: 2f97 al driver destino [2][5], en modo 1
UVM_INFO Driver.sv(59) @ 1110: uvm_test_top.amb_inst.agent.drv_inst11 [DRV] Driver #11: Fuente: [5][4], envia el mensaje: 1f92 al driver destino [5][4], en modo 1

UVM_INFO monitor.sv(40) @ 550: uvm_test_top.amb_inst.agent.mnt_inst15 [Monitor] Monitor #15: Destino: [4][5] recibe dato: 3a5d de drvr fuente [4][5] en modo 1
UVM_INFO monitor.sv(40) @ 630: uvm_test_top.amb_inst.agent.mnt_inst9 [Monitor] Monitor #9: Destino: [5][2] recibe dato: 3500 de drvr fuente [0][2] en modo 0
UVM_INFO monitor.sv(40) @ 790: uvm_test_top.amb_inst.agent.mnt_inst14 [Monitor] Monitor #14: Destino: [3][5] recibe dato: 441c de drvr fuente [4][0] en modo 1
UVM_INFO monitor.sv(40) @ 1110: uvm_test_top.amb_inst.agent.mnt_inst10 [Monitor] Monitor #10: Destino: [5][3] recibe dato: 1d35 de drvr fuente [0][4] en modo 1
UVM_INFO monitor.sv(40) @ 1150: uvm_test_top.amb_inst.agent.mnt_inst11 [Monitor] Monitor #11: Destino: [5][4] recibe dato: 1f92 de drvr fuente [5][4] en modo 1
UVM_INFO monitor.sv(40) @ 1230: uvm_test_top.amb_inst.agent.mnt_inst10 [Monitor] Monitor #10: Destino: [5][3] recibe dato: 2a94 de drvr fuente [3][0] en modo 1
UVM_INFO monitor.sv(40) @ 1270: uvm_test_top.amb_inst.agent.mnt_inst11 [Monitor] Monitor #11: Destino: [5][4] recibe dato: 518d de drvr fuente [3][5] en modo 1
UVM_INFO monitor.sv(40) @ 1910: uvm_test_top.amb_inst.agent.mnt_inst12 [Monitor] Monitor #12: Destino: [1][5] recibe dato: 6fcf de drvr fuente [2][0] en modo 0*/