class Item extends uvm_sequence_item;

    `uvm_object_utils(Item);

    function new(string name = "Item");
    